`timescale 1ns / 1ps

module tb_adder();

    reg a3,a2,a1,a0,b3,b2,b1,b0,cin;//input
    wire s3,s2,s1,s0, cout;//output

fb_adder duts(
    .a3(a3),
    .a2(a2),
    .a1(a1),
    .a0(a0),
    .b3(b3),
    .b2(b2),
    .b1(b1),
    .b0(b0),
    .cin(cin),
    .s3(s3),
    .s2(s2),
    .s1(s1),
    .s0(s0),
    .cout(cout)
);

initial begin
    
    #0;
    a3 = 1'b0; a2 = 1'b0; a1 = 1'b0; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    cin = 1'b0;
    #1;//delay 값 유지
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b0; a1 = 1'b0; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b0; a1 = 1'b1; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b0; a1 = 1'b1; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b0; a0 = 1'b0;   
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b0; a0 = 1'b1;  
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b1; a0 = 1'b0;  
     b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b1; a0 = 1'b1;  
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b0; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b0; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b1; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b1; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b1; a1 = 1'b0; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b1; a1 = 1'b1; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b1; a1 = 1'b1; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    $finish;
end

endmodule
